
interface intf();
    // ------------------- port declaration-------------------------------------
    logic [3:0]  in;
    logic [6:0] out;
    //--------------------------------------------------------------------------
endinterface

